library verilog;
use verilog.vl_types.all;
entity topLevel_vlg_vec_tst is
end topLevel_vlg_vec_tst;
